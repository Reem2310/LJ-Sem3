<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-53.927,-20.7762,98.5273,-96.1315</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>17.5,-47.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>16.5,-40.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_INVERTER</type>
<position>-94.5,-27.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,-48.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-39.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-41.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>25,-40.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>25,-47.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>12,-35.5</position>
<gparam>LABEL_TEXT Half-Substractor(2-input 1-bit)</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-60.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>2.5,-60.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>9.5,-60.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>20,-67</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>20,-72.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>20,-78</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_OR3</type>
<position>33,-72.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR3</type>
<position>20.5,-86</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>10 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1.5,-66</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_INVERTER</type>
<position>-102,-47</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>42,-72.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>31,-86</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>11.5,-56</position>
<gparam>LABEL_TEXT Full-Subtractor(3-input 1-bit))</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-39.5,13.5,-39.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>5.5 2</intersection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5.5,-48.5,5.5,-39.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-39.5,13.5,-39.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-41.5,13.5,-41.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>8 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,-46.5,8,-41.5</points>
<intersection>-46.5 5</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>8,-46.5,14.5,-46.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>8 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-48.5,14.5,-48.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-47.5,24,-47.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-40.5,24,-40.5</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,-66,17,-66</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>1.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>1.5,-71.5,1.5,-66</points>
<intersection>-71.5 7</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>1.5,-71.5,17,-71.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>1.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-86,2.5,-62.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-86 5</intersection>
<intersection>-77 3</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-68,17,-68</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-77,17,-77</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>2.5,-86,17.5,-86</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-88,9.5,-62.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-88 5</intersection>
<intersection>-79 3</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-73.5,17,-73.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>9.5,-79,17,-79</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>9.5,-88,17.5,-88</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-84,-4.5,-62.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-84 3</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-66,-3.5,-66</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-84,17.5,-84</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-70.5,26.5,-67</points>
<intersection>-70.5 1</intersection>
<intersection>-67 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-70.5,30,-70.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-67,26.5,-67</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-72.5,30,-72.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-78,26.5,-74.5</points>
<intersection>-78 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-78,26.5,-78</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-74.5,30,-74.5</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-72.5,41,-72.5</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-86,30,-86</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>34</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>