<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-473.171,171.715,-333.907,97.5875</PageViewport>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>-411,106</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-421.5,106</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>-400,106</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-412,113</position>
<gparam>LABEL_TEXT All Gate's Using Universal Gate NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>-430.5,106.5</position>
<gparam>LABEL_TEXT NOT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>-411,97.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>-395.5,97.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>-421.5,97.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>-385,97.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>-430.5,98</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>BA_NAND2</type>
<position>-411,88</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>-411,82.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>BA_NAND2</type>
<position>-398.5,85.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-421.5,88</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-421.5,82.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>-387.5,85.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>-430.5,86.5</position>
<gparam>LABEL_TEXT OR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>-411,74.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>BA_NAND2</type>
<position>-411,67.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>BA_NAND2</type>
<position>-398.5,71.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND2</type>
<position>-386,71.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>-421.5,74.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>-421.5,67.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>-376,71.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>-430,72</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>BA_NAND2</type>
<position>-411,59.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>BA_NAND2</type>
<position>-411,45.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>BA_NAND2</type>
<position>-398,54</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>-397.5,36</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>-383,48</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>-423.5,52</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>-423.5,46.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>-372.5,48</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>-430.5,49.5</position>
<gparam>LABEL_TEXT EX-OR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>-411,24</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>-410.5,10</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>-394.5,19</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BA_NAND2</type>
<position>-401,3</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_NAND2</type>
<position>-380.5,12</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>-429.5,25</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>-429.5,11</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>-369,12</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-437.5,16</position>
<gparam>LABEL_TEXT EX-NOR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,105,-416.5,107</points>
<intersection>105 4</intersection>
<intersection>106 2</intersection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,107,-414,107</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-419.5,106,-416.5,106</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-416.5,105,-414,105</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-408,106,-401,106</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,96.5,-416.5,98.5</points>
<intersection>96.5 4</intersection>
<intersection>97.5 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,98.5,-414,98.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-419.5,97.5,-416.5,97.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-416.5,96.5,-414,96.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,96.5,-403,98.5</points>
<intersection>96.5 4</intersection>
<intersection>97.5 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403,98.5,-398.5,98.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,97.5,-403,97.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-403 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-403,96.5,-398.5,96.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-403 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-392.5,97.5,-386,97.5</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,87,-416.5,89</points>
<intersection>87 1</intersection>
<intersection>88 2</intersection>
<intersection>89 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,87,-414,87</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-419.5,88,-416.5,88</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-416.5,89,-414,89</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,81.5,-416.5,83.5</points>
<intersection>81.5 5</intersection>
<intersection>82.5 1</intersection>
<intersection>83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-419.5,82.5,-416.5,82.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-416.5,83.5,-414,83.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-416.5,81.5,-414,81.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404.5,86.5,-404.5,88</points>
<intersection>86.5 1</intersection>
<intersection>88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-404.5,86.5,-401.5,86.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-404.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,88,-404.5,88</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>-404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404.5,82.5,-404.5,84.5</points>
<intersection>82.5 1</intersection>
<intersection>84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-408,82.5,-404.5,82.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-404.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-404.5,84.5,-401.5,84.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-395.5,85.5,-388.5,85.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,73.5,-416.5,75.5</points>
<intersection>73.5 4</intersection>
<intersection>74.5 2</intersection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,75.5,-414,75.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-419.5,74.5,-416.5,74.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-416.5,73.5,-414,73.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,66.5,-416.5,68.5</points>
<intersection>66.5 4</intersection>
<intersection>67.5 2</intersection>
<intersection>68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,68.5,-414,68.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-419.5,67.5,-416.5,67.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-416.5,66.5,-414,66.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404.5,72.5,-404.5,74.5</points>
<intersection>72.5 1</intersection>
<intersection>74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-404.5,72.5,-401.5,72.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-404.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,74.5,-404.5,74.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>-404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404.5,67.5,-404.5,70.5</points>
<intersection>67.5 1</intersection>
<intersection>70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-408,67.5,-404.5,67.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>-404.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-404.5,70.5,-401.5,70.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-404.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-392,70.5,-392,72.5</points>
<intersection>70.5 4</intersection>
<intersection>71.5 2</intersection>
<intersection>72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-392,72.5,-389,72.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-392 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395.5,71.5,-392,71.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>-392 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-392,70.5,-389,70.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-392 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-383,71.5,-377,71.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>44</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-417.5,35,-417.5,60.5</points>
<intersection>35 6</intersection>
<intersection>52 2</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-417.5,60.5,-414,60.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-417.5 0</intersection>
<intersection>-414 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-421.5,52,-417.5,52</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-417.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-417.5,35,-400.5,35</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-417.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-414,58.5,-414,60.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>60.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-401,55,-401,59.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>59.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-408,59.5,-401,59.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-401 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404,37,-404,45.5</points>
<intersection>37 1</intersection>
<intersection>45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-404,37,-400.5,37</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-404 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,45.5,-404,45.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-404 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-390,36,-390,47</points>
<intersection>36 2</intersection>
<intersection>47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-390,47,-386,47</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-390 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-394.5,36,-390,36</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-390 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-390.5,49,-390.5,54</points>
<intersection>49 1</intersection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-390.5,49,-386,49</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-390.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395,54,-390.5,54</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>-390.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-380,48,-373.5,48</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-415.5,44.5,-415.5,53</points>
<intersection>44.5 1</intersection>
<intersection>53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-415.5,44.5,-414,44.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-415.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-415.5,53,-401,53</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-415.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-421.5,46.5,-414,46.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-427.5,25,-414,25</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-425.5 3</intersection>
<intersection>-414 10</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-425.5,2,-425.5,25</points>
<intersection>2 6</intersection>
<intersection>25 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-425.5,2,-404,2</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>-425.5 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-414,23,-414,25</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>25 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-417,9,-417,18</points>
<intersection>9 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-417,18,-397.5,18</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-417 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-417,9,-413.5,9</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-417 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-402.5,20,-402.5,24</points>
<intersection>20 1</intersection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-402.5,20,-397.5,20</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,24,-402.5,24</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-427.5,11,-413.5,11</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-405.5,4,-405.5,10</points>
<intersection>4 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-405.5,4,-404,4</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-405.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-407.5,10,-405.5,10</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-387.5,13,-387.5,19</points>
<intersection>13 1</intersection>
<intersection>19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-387.5,13,-383.5,13</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-387.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-391.5,19,-387.5,19</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>-387.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-390.5,3,-390.5,11</points>
<intersection>3 2</intersection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-390.5,11,-383.5,11</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>-390.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-398,3,-390.5,3</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>-390.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-377.5,12,-370,12</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<connection>
<GID>80</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-11.6485,91.3706,127.458,17.3267</PageViewport>
<gate>
<ID>90</ID>
<type>BE_NOR2</type>
<position>42,69.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>31.5,69.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>52,69.5</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>24,69.5</position>
<gparam>LABEL_TEXT NOT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>38.5,78</position>
<gparam>LABEL_TEXT ALL Gate's Using NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>100</ID>
<type>BE_NOR2</type>
<position>42,60.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>BE_NOR2</type>
<position>42,53</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>BE_NOR2</type>
<position>53.5,57</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>31.5,60.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>31.5,53</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>63,57</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>24,58</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>BE_NOR2</type>
<position>42,45</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>BE_NOR2</type>
<position>54,45</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>31.5,45</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>65,45</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>24.5,45</position>
<gparam>LABEL_TEXT OR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>BE_NOR2</type>
<position>42,34.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>BE_NOR2</type>
<position>42,26</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>BE_NOR2</type>
<position>52.5,30.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>BE_NOR2</type>
<position>66.5,30.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>31.5,34.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>31.5,26</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>75,30.5</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>24,30.5</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>BE_NOR2</type>
<position>41.5,14</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>BE_NOR2</type>
<position>71,13</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>BE_NOR2</type>
<position>83.5,7</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>100.5,7</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>BE_NOR2</type>
<position>42,-7.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>BE_NOR2</type>
<position>59,-1</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>30,14</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>30.5,-8.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>111,7</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>23.5,4</position>
<gparam>LABEL_TEXT XOR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BE_NOR2</type>
<position>54,-26.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>BE_NOR2</type>
<position>54,-36</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>BE_NOR2</type>
<position>54,-46</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>BE_NOR2</type>
<position>69,-41</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>BE_NOR2</type>
<position>84.5,-35.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>BE_NOR2</type>
<position>101,-35.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>33.5,-25.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_TOGGLE</type>
<position>38.5,-30</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>113,-35.5</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>24,-34</position>
<gparam>LABEL_TEXT X-NOR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,68.5,36,70.5</points>
<intersection>68.5 4</intersection>
<intersection>69.5 2</intersection>
<intersection>70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,70.5,39,70.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,69.5,36,69.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,68.5,39,68.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,69.5,51,69.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,59.5,36,61.5</points>
<intersection>59.5 4</intersection>
<intersection>60.5 2</intersection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,61.5,39,61.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,60.5,36,60.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,59.5,39,59.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,52,36,54</points>
<intersection>52 4</intersection>
<intersection>53 2</intersection>
<intersection>54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,54,39,54</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,53,36,53</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,52,39,52</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,58,47.5,60.5</points>
<intersection>58 1</intersection>
<intersection>60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,58,50.5,58</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,60.5,47.5,60.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,53,47.5,56</points>
<intersection>53 1</intersection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,53,47.5,53</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,56,50.5,56</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,57,62,57</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,44,36,46</points>
<intersection>44 4</intersection>
<intersection>45 2</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,46,39,46</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,45,36,45</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,44,39,44</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,44,48,46</points>
<intersection>44 4</intersection>
<intersection>45 2</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,46,51,46</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,45,48,45</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>48,44,51,44</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,45,64,45</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>120</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,33.5,36,35.5</points>
<intersection>33.5 4</intersection>
<intersection>34.5 2</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,35.5,39,35.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,34.5,36,34.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,33.5,39,33.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,25,36,27</points>
<intersection>25 4</intersection>
<intersection>26 2</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,27,39,27</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,26,36,26</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,25,39,25</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,31.5,47,34.5</points>
<intersection>31.5 1</intersection>
<intersection>34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,31.5,49.5,31.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,34.5,47,34.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,26,47,29.5</points>
<intersection>26 1</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,26,47,26</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,29.5,49.5,29.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,29.5,59.5,31.5</points>
<intersection>29.5 4</intersection>
<intersection>30.5 2</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,31.5,63.5,31.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,30.5,59.5,30.5</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>59.5,29.5,63.5,29.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,30.5,74,30.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<connection>
<GID>136</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,7,110,7</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>156</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,0,38.5,15</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>0 6</intersection>
<intersection>14 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>38.5,0,56,0</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>32,14,38.5,14</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-10.5,35.5,-8.5</points>
<intersection>-10.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-10.5,68,-10.5</points>
<intersection>35.5 0</intersection>
<intersection>39 6</intersection>
<intersection>68 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-8.5,39,-8.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection>
<intersection>39 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>68,-10.5,68,12</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>39,-10.5,39,-6.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-7.5,50.5,-2</points>
<intersection>-7.5 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-2,56,-2</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-7.5,50.5,-7.5</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,14,68,14</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,8,77,13</points>
<intersection>8 1</intersection>
<intersection>13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,8,80.5,8</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,13,77,13</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-1,71,6</points>
<intersection>-1 1</intersection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-1,71,-1</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,6,80.5,6</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,6,92,8</points>
<intersection>6 4</intersection>
<intersection>7 2</intersection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,8,97.5,8</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,7,92,7</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>92,6,97.5,6</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-25.5,51,-25.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>35.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>35.5,-46,35.5,-25.5</points>
<intersection>-46 3</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>35.5,-46,51,-46</points>
<intersection>35.5 2</intersection>
<intersection>51 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51,-47,51,-45</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-46 3</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-36,45,-27.5</points>
<intersection>-36 4</intersection>
<intersection>-30 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-27.5,51,-27.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-30,45,-30</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>45,-36,51,-36</points>
<intersection>45 0</intersection>
<intersection>51 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>51,-37,51,-35</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-36 4</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-34.5,69,-26.5</points>
<intersection>-34.5 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-34.5,81.5,-34.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-26.5,69,-26.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-41,76.5,-36.5</points>
<intersection>-41 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-36.5,81.5,-36.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-41,76.5,-41</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-40,61.5,-36</points>
<intersection>-40 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61.5,-40,66,-40</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-36,61.5,-36</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-46,61.5,-42</points>
<intersection>-46 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-46,61.5,-46</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-42,66,-42</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-36.5,92.5,-34.5</points>
<intersection>-36.5 4</intersection>
<intersection>-35.5 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-34.5,98,-34.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-35.5,92.5,-35.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>92.5,-36.5,98,-36.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-35.5,112,-35.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>176</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-477.177,289.746,916.823,-452.254</PageViewport></page 2>
<page 3>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 3>
<page 4>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 4>
<page 5>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 5>
<page 6>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 6>
<page 7>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 7>
<page 8>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 8>
<page 9>
<PageViewport>0,35.7538,439.646,-198.262</PageViewport></page 9></circuit>