<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-45.7875,-25.927,81.0125,-88.6019</PageViewport>
<gate>
<ID>2</ID>
<type>AI_XOR2</type>
<position>3,-51.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>26.5,-52.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>8.5,-63</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-50.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-52.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-68.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>28.5,-63.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR2</type>
<position>44.5,-70</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>52,-52.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>52,-70</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>16.5,-43</position>
<gparam>LABEL_TEXT Alternative Equation Half Using of Full-Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-50.5,0,-50.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-64,-6,-50.5</points>
<intersection>-64 4</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-6,-64,5.5,-64</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-6 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-52.5,0,-52.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-62,-1.5,-52.5</points>
<intersection>-62 4</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-1.5,-62,5.5,-62</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-1.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-51.5,23.5,-51.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-62.5,18,-51.5</points>
<intersection>-62.5 4</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>18,-62.5,25.5,-62.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>18 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-71,13.5,-63</points>
<intersection>-71 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-71,41.5,-71</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-63,13.5,-63</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-69,36.5,-63.5</points>
<intersection>-69 1</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-69,41.5,-69</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-63.5,36.5,-63.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-68.5,21,-53.5</points>
<intersection>-68.5 2</intersection>
<intersection>-64.5 3</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-53.5,23.5,-53.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-68.5,21,-68.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21,-64.5,25.5,-64.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-70,51,-70</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-52.5,51,-52.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>