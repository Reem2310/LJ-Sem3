<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-24.0326,-25.927,102.767,-88.6019</PageViewport>
<gate>
<ID>2</ID>
<type>AI_XOR2</type>
<position>6.5,-52</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>28,-53</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>7,-66.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>31.5,-69.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>46,-75.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-4,-51</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-4,-53</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-3.5,-74.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>1,-65.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>24.5,-68.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>38.5,-53</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>53,-75.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>17.5,-44</position>
<gparam>LABEL_TEXT Alternate Equation (FS Using HS)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-51,3.5,-51</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-1 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1,-65.5,-1,-51</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-53,3.5,-53</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-2 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-2,-67.5,-2,-53</points>
<intersection>-67.5 4</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-2,-67.5,4,-67.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-2 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-65.5,4,-65.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-74.5,20,-54</points>
<intersection>-74.5 1</intersection>
<intersection>-70.5 3</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-74.5,20,-74.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-54,25,-54</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>20,-70.5,28.5,-70.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-76.5,15,-66.5</points>
<intersection>-76.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-76.5,43,-76.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-66.5,15,-66.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26.5,-68.5,28.5,-68.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-52,25,-52</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-68.5,17,-52</points>
<intersection>-68.5 4</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-68.5,22.5,-68.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>17 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-74.5,38.5,-69.5</points>
<intersection>-74.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-74.5,43,-74.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-69.5,38.5,-69.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-75.5,52,-75.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-53,37.5,-53</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>